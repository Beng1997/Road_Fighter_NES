

 module menu_textBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output	logic	[3:0] HitEdgeCode //one bit per edge 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] COLOR_ENCODING = 8'hFF ;// RGB value in the bitmap representing the BITMAP coolor
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:63][0:255] object_colors = {
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111000000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111000000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111000000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111000000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111000000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110001111111111100000000000011111111101111111111110000111111100011111111111000001111111111111,
	256'b1111111111000011111111111000001111111111110000111111111000011111111100000001111111111110111111000001101111111111111011111111111110111111111110000000000011111111111110111111111111111000000000011111111101111111111110011111111111011111111111000001111111111111,
	256'b1110000000110011000000000111001100000000000011000000000011100000000000000001100000000000111111000001100000011100000011100000000000110000000001110000000000000111000000111000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111111000001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111111000001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111111000001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111111000001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111000110001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111000110001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111000110001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000110001100000000000011000000000011100000000000000001100000000000111000110001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1110000000110011000000000111001100000000000011000000000011100000000000000001100000000000111000110001100000011100000011100000000000110000000001110000000000000111000000110000000000111000000011100000000000000011100000011000000111011100000000111000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000110001100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000001111100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000001111100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000001111100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000001111100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1111111111000011111111111000001111110000000000111111100000011111100000000001111110000000111000001111100000011100000011111100000000111111111110000000000000000111000000110000000000111000000000011111100000000011100000011111111111011111111111000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000001111100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000001111100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000001111100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000001111100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000001111100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000001110000001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000011100000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000110000000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000110000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000001100001100000000000000000000111000000000011100000001100000000000111000000001100000011100000011100000000000110000000011000000000000000111000000111000000000111000000000000000011100000011100000011000000111011100000001110000000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000,
	256'b1110000000000011000000000011101111111111110011111111100011111111100000000001111111111110111000000001100000011100000011111111111110110000000000111000000000000111000000001111111111100000000011111111100000000011100000011000000111011100000000001100000011100000};

 
 
//////////--------------------------------------------------------------------------------------------------------------= 
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
//there is one bit per edge, in the corner two bits are set  
 logic [0:3] [0:3] [3:0] hit_colors = 
		   {16'hC446,     
			16'h8C62,    
			16'h8932, 
			16'h9113}; 
 // pipeline (ff) to get the pixel color from the array 	 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) begin 
		RGBout <=	8'h00; 
		HitEdgeCode <= 4'h0; 
	end 
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default  
		HitEdgeCode <= 4'h0; 
 
		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket  
			HitEdgeCode <= hit_colors[offsetY >> 4][offsetX >> 6 ]; // get hitting edge from the colors table
			RGBout <= (object_colors[offsetY][offsetX] ==  1 ) ? COLOR_ENCODING  : TRANSPARENT_ENCODING; 
		end  	 
		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
