
 module winBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY, 
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
 
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output	logic	[3:0] HitEdgeCode //one bit per edge 
 ) ; 
 
 
// generating the bitmap 
 

localparam logic [7:0] COLOR_ENCODING = 8'hFF ;// RGB value in the bitmap representing the BITMAP coolor
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:63][0:127] object_colors = {
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111100000000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111100000000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111100000000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111100000000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111100000000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b11100000000000111100000111111111111111000000011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b11100000000000111100111111111111111111111100011110000000001111000000000001110000000000011110000111111100111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111111100000001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00011110000111000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100011110001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000000000011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000001111111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001110000111100011110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111001110,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111000000,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111000000,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111000000,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111000000,
	128'b00000001111000000000111000000000000000111100011110000000001111000000000001111111000011111110000011110000111100000000001111000000,
	128'b00000001111000000000000011111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110,
	128'b00000001111000000000000111111111111111000000000001111111110000000000000001110000000000011110000111111100111100000000001111001110};

 
 
//////////--------------------------------------------------------------------------------------------------------------= 
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
//there is one bit per edge, in the corner two bits are set  
 logic [0:3] [0:3] [3:0] hit_colors = 
		   {16'hC446,     
			16'h8C62,    
			16'h8932, 
			16'h9113}; 
 // pipeline (ff) to get the pixel color from the array 	 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) begin 
		RGBout <=	8'h00; 
		HitEdgeCode <= 4'h0; 
	end 
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default  
		HitEdgeCode <= 4'h0; 
 
		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket  
			HitEdgeCode <= hit_colors[offsetY >> 4][offsetX >> 5 ]; // get hitting edge from the colors table
			RGBout <= (object_colors[offsetY][offsetX] ==  1 ) ? COLOR_ENCODING  : TRANSPARENT_ENCODING; 
		end  	 
		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
